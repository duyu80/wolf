//************************************************************************
//**                          Baseboard CPLD							**
//**                          PRSNT_LED_CTRL.v						    **
//************************************************************************ 

//**********************      ChangeList      *****************************

`include "../SRC/baseboard_define.v"

module PRSNT_LED_CTRL (
            // System
			input      SYSCLK,
			input      RESET_N,
            // Driver present and amber LED inout
			inout      DRV3_PRSNT_AMBER_LED,DRV2_PRSNT_AMBER_LED,DRV1_PRSNT_AMBER_LED,DRV0_PRSNT_AMBER_LED,
			inout      DRV7_PRSNT_AMBER_LED,DRV6_PRSNT_AMBER_LED,DRV5_PRSNT_AMBER_LED,DRV4_PRSNT_AMBER_LED,
			inout      DRV11_PRSNT_AMBER_LED,DRV10_PRSNT_AMBER_LED,DRV9_PRSNT_AMBER_LED,DRV8_PRSNT_AMBER_LED,
			inout      DRV15_PRSNT_AMBER_LED,DRV14_PRSNT_AMBER_LED,DRV13_PRSNT_AMBER_LED,DRV12_PRSNT_AMBER_LED,
			inout      DRV19_PRSNT_AMBER_LED,DRV18_PRSNT_AMBER_LED,DRV17_PRSNT_AMBER_LED,DRV16_PRSNT_AMBER_LED,
			inout      DRV23_PRSNT_AMBER_LED,DRV22_PRSNT_AMBER_LED,DRV21_PRSNT_AMBER_LED,DRV20_PRSNT_AMBER_LED,
			inout      DRV27_PRSNT_AMBER_LED,DRV26_PRSNT_AMBER_LED,DRV25_PRSNT_AMBER_LED,DRV24_PRSNT_AMBER_LED,
			inout      DRV31_PRSNT_AMBER_LED,DRV30_PRSNT_AMBER_LED,DRV29_PRSNT_AMBER_LED,DRV28_PRSNT_AMBER_LED,
			inout      DRV35_PRSNT_AMBER_LED,DRV34_PRSNT_AMBER_LED,DRV33_PRSNT_AMBER_LED,DRV32_PRSNT_AMBER_LED,
            // Driver identify and blue LED inout
			inout      DRV3_IFDET_BLUE_LED,DRV2_IFDET_BLUE_LED,DRV1_IFDET_BLUE_LED,DRV0_IFDET_BLUE_LED,
			inout      DRV7_IFDET_BLUE_LED,DRV6_IFDET_BLUE_LED,DRV5_IFDET_BLUE_LED,DRV4_IFDET_BLUE_LED,
			inout      DRV11_IFDET_BLUE_LED,DRV10_IFDET_BLUE_LED,DRV9_IFDET_BLUE_LED,DRV8_IFDET_BLUE_LED,
			inout      DRV15_IFDET_BLUE_LED,DRV14_IFDET_BLUE_LED,DRV13_IFDET_BLUE_LED,DRV12_IFDET_BLUE_LED,
			inout      DRV19_IFDET_BLUE_LED,DRV18_IFDET_BLUE_LED,DRV17_IFDET_BLUE_LED,DRV16_IFDET_BLUE_LED,
			inout      DRV23_IFDET_BLUE_LED,DRV22_IFDET_BLUE_LED,DRV21_IFDET_BLUE_LED,DRV20_IFDET_BLUE_LED,
			inout      DRV27_IFDET_BLUE_LED,DRV26_IFDET_BLUE_LED,DRV25_IFDET_BLUE_LED,DRV24_IFDET_BLUE_LED,
			inout      DRV31_IFDET_BLUE_LED,DRV30_IFDET_BLUE_LED,DRV29_IFDET_BLUE_LED,DRV28_IFDET_BLUE_LED,
			inout      DRV35_IFDET_BLUE_LED,DRV34_IFDET_BLUE_LED,DRV33_IFDET_BLUE_LED,DRV32_IFDET_BLUE_LED,
            // Amber LED data
			input      [35:0]    AMBER_DAT,
            // Blue LED data
            input      [35:0]    BLUE_DAT,			
            // Present signal
			output reg [35:0]    PRSNT,
			// Identify signal
			output reg [35:0]    IDENT
			);

reg    [31:0]  CNT;
reg    [35:0]  DRV_PRSNT_AMBER_LED_EN;
reg    [35:0]  DRV_IFDET_BLUE_LED_EN;

always@(posedge SYSCLK or negedge RESET_N)
	begin
		if(RESET_N == 1'b0)
			begin
			    CNT                    <= 32'h0;
				DRV_PRSNT_AMBER_LED_EN <= 36'h0;
				DRV_IFDET_BLUE_LED_EN  <= 36'h0;
			end
		else
		    begin
			    CNT                    <= (CNT < `TIME_100MS)? (CNT + 32'd1) : 32'd0;
				DRV_PRSNT_AMBER_LED_EN <= (CNT < `TIME_99MS)? 36'hf_ffff_ffff : 36'h0;
				DRV_IFDET_BLUE_LED_EN  <= (CNT < `TIME_99MS)? 36'hf_ffff_ffff : 36'h0;
			end
	end

always@(posedge SYSCLK or negedge RESET_N)
	begin
		if(RESET_N == 1'b0)
			begin
			    PRSNT <= 36'h0;
				IDENT <= 36'h0;
			end
		else
		    begin
			
			    PRSNT <= (CNT == `TIME_100MS)? {
			    ~DRV35_IFDET_BLUE_LED,~DRV34_IFDET_BLUE_LED,~DRV33_IFDET_BLUE_LED,~DRV32_IFDET_BLUE_LED,			
			    ~DRV31_IFDET_BLUE_LED,~DRV30_IFDET_BLUE_LED,~DRV29_IFDET_BLUE_LED,~DRV28_IFDET_BLUE_LED,			
			    ~DRV27_IFDET_BLUE_LED,~DRV26_IFDET_BLUE_LED,~DRV25_IFDET_BLUE_LED,~DRV24_IFDET_BLUE_LED,			
			    ~DRV23_IFDET_BLUE_LED,~DRV22_IFDET_BLUE_LED,~DRV21_IFDET_BLUE_LED,~DRV20_IFDET_BLUE_LED,			
			    ~DRV19_IFDET_BLUE_LED,~DRV18_IFDET_BLUE_LED,~DRV17_IFDET_BLUE_LED,~DRV16_IFDET_BLUE_LED,			
			    ~DRV15_IFDET_BLUE_LED,~DRV14_IFDET_BLUE_LED,~DRV13_IFDET_BLUE_LED,~DRV12_IFDET_BLUE_LED,			
			    ~DRV11_IFDET_BLUE_LED,~DRV10_IFDET_BLUE_LED,~DRV9_IFDET_BLUE_LED,~DRV8_IFDET_BLUE_LED,			
			    ~DRV7_IFDET_BLUE_LED,~DRV6_IFDET_BLUE_LED,~DRV5_IFDET_BLUE_LED,~DRV4_IFDET_BLUE_LED,			
                ~DRV3_IFDET_BLUE_LED,~DRV2_IFDET_BLUE_LED,~DRV1_IFDET_BLUE_LED,~DRV0_IFDET_BLUE_LED
                } : PRSNT;
				
                IDENT <= (CNT == `TIME_100MS)? {
			    DRV35_PRSNT_AMBER_LED,DRV34_PRSNT_AMBER_LED,DRV33_PRSNT_AMBER_LED,DRV32_PRSNT_AMBER_LED,			
			    DRV31_PRSNT_AMBER_LED,DRV30_PRSNT_AMBER_LED,DRV29_PRSNT_AMBER_LED,DRV28_PRSNT_AMBER_LED,			
			    DRV27_PRSNT_AMBER_LED,DRV26_PRSNT_AMBER_LED,DRV25_PRSNT_AMBER_LED,DRV24_PRSNT_AMBER_LED,			
			    DRV23_PRSNT_AMBER_LED,DRV22_PRSNT_AMBER_LED,DRV21_PRSNT_AMBER_LED,DRV20_PRSNT_AMBER_LED,			
			    DRV19_PRSNT_AMBER_LED,DRV18_PRSNT_AMBER_LED,DRV17_PRSNT_AMBER_LED,DRV16_PRSNT_AMBER_LED,			
			    DRV15_PRSNT_AMBER_LED,DRV14_PRSNT_AMBER_LED,DRV13_PRSNT_AMBER_LED,DRV12_PRSNT_AMBER_LED,			
			    DRV11_PRSNT_AMBER_LED,DRV10_PRSNT_AMBER_LED,DRV9_PRSNT_AMBER_LED,DRV8_PRSNT_AMBER_LED,			
			    DRV7_PRSNT_AMBER_LED,DRV6_PRSNT_AMBER_LED,DRV5_PRSNT_AMBER_LED,DRV4_PRSNT_AMBER_LED,			
                DRV3_PRSNT_AMBER_LED,DRV2_PRSNT_AMBER_LED,DRV1_PRSNT_AMBER_LED,DRV0_PRSNT_AMBER_LED
                } : IDENT;

			end
	end


assign    DRV0_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[0]? AMBER_DAT[0] : 1'bz;
assign    DRV1_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[1]? AMBER_DAT[1] : 1'bz;
assign    DRV2_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[2]? AMBER_DAT[2] : 1'bz;
assign    DRV3_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[3]? AMBER_DAT[3] : 1'bz;
assign    DRV4_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[4]? AMBER_DAT[4] : 1'bz;
assign    DRV5_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[5]? AMBER_DAT[5] : 1'bz;
assign    DRV6_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[6]? AMBER_DAT[6] : 1'bz;
assign    DRV7_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[7]? AMBER_DAT[7] : 1'bz;
assign    DRV8_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[8]? AMBER_DAT[8] : 1'bz;
assign    DRV9_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[9]? AMBER_DAT[9] : 1'bz;
assign    DRV10_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[10]? AMBER_DAT[10] : 1'bz;
assign    DRV11_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[11]? AMBER_DAT[11] : 1'bz;
assign    DRV12_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[12]? AMBER_DAT[12] : 1'bz;
assign    DRV13_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[13]? AMBER_DAT[13] : 1'bz;
assign    DRV14_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[14]? AMBER_DAT[14] : 1'bz;
assign    DRV15_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[15]? AMBER_DAT[15] : 1'bz;
assign    DRV16_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[16]? AMBER_DAT[16] : 1'bz;
assign    DRV17_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[17]? AMBER_DAT[17] : 1'bz;
assign    DRV18_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[18]? AMBER_DAT[18] : 1'bz;
assign    DRV19_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[19]? AMBER_DAT[19] : 1'bz;
assign    DRV20_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[20]? AMBER_DAT[20] : 1'bz;
assign    DRV21_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[21]? AMBER_DAT[21] : 1'bz;
assign    DRV22_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[22]? AMBER_DAT[22] : 1'bz;
assign    DRV23_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[23]? AMBER_DAT[23] : 1'bz;
assign    DRV24_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[24]? AMBER_DAT[24] : 1'bz;
assign    DRV25_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[25]? AMBER_DAT[25] : 1'bz;
assign    DRV26_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[26]? AMBER_DAT[26] : 1'bz;
assign    DRV27_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[27]? AMBER_DAT[27] : 1'bz;
assign    DRV28_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[28]? AMBER_DAT[28] : 1'bz;
assign    DRV29_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[29]? AMBER_DAT[29] : 1'bz;
assign    DRV30_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[30]? AMBER_DAT[30] : 1'bz;
assign    DRV31_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[31]? AMBER_DAT[31] : 1'bz;
assign    DRV32_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[32]? AMBER_DAT[32] : 1'bz;
assign    DRV33_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[33]? AMBER_DAT[33] : 1'bz;
assign    DRV34_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[34]? AMBER_DAT[34] : 1'bz;
assign    DRV35_PRSNT_AMBER_LED = DRV_PRSNT_AMBER_LED_EN[35]? AMBER_DAT[35] : 1'bz;

assign    DRV0_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[0]? BLUE_DAT[0] : 1'bz;
assign    DRV1_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[1]? BLUE_DAT[1] : 1'bz;
assign    DRV2_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[2]? BLUE_DAT[2] : 1'bz;
assign    DRV3_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[3]? BLUE_DAT[3] : 1'bz;
assign    DRV4_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[4]? BLUE_DAT[4] : 1'bz;
assign    DRV5_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[5]? BLUE_DAT[5] : 1'bz;
assign    DRV6_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[6]? BLUE_DAT[6] : 1'bz;
assign    DRV7_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[7]? BLUE_DAT[7] : 1'bz;
assign    DRV8_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[8]? BLUE_DAT[8] : 1'bz;
assign    DRV9_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[9]? BLUE_DAT[9] : 1'bz;
assign    DRV10_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[10]? BLUE_DAT[10] : 1'bz;
assign    DRV11_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[11]? BLUE_DAT[11] : 1'bz;
assign    DRV12_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[12]? BLUE_DAT[12] : 1'bz;
assign    DRV13_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[13]? BLUE_DAT[13] : 1'bz;
assign    DRV14_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[14]? BLUE_DAT[14] : 1'bz;
assign    DRV15_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[15]? BLUE_DAT[15] : 1'bz;
assign    DRV16_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[16]? BLUE_DAT[16] : 1'bz;
assign    DRV17_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[17]? BLUE_DAT[17] : 1'bz;
assign    DRV18_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[18]? BLUE_DAT[18] : 1'bz;
assign    DRV19_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[19]? BLUE_DAT[19] : 1'bz;
assign    DRV20_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[20]? BLUE_DAT[20] : 1'bz;
assign    DRV21_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[21]? BLUE_DAT[21] : 1'bz;
assign    DRV22_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[22]? BLUE_DAT[22] : 1'bz;
assign    DRV23_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[23]? BLUE_DAT[23] : 1'bz;
assign    DRV24_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[24]? BLUE_DAT[24] : 1'bz;
assign    DRV25_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[25]? BLUE_DAT[25] : 1'bz;
assign    DRV26_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[26]? BLUE_DAT[26] : 1'bz;
assign    DRV27_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[27]? BLUE_DAT[27] : 1'bz;
assign    DRV28_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[28]? BLUE_DAT[28] : 1'bz;
assign    DRV29_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[29]? BLUE_DAT[29] : 1'bz;
assign    DRV30_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[30]? BLUE_DAT[30] : 1'bz;
assign    DRV31_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[31]? BLUE_DAT[31] : 1'bz;
assign    DRV32_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[32]? BLUE_DAT[32] : 1'bz;
assign    DRV33_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[33]? BLUE_DAT[33] : 1'bz;
assign    DRV34_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[34]? BLUE_DAT[34] : 1'bz;
assign    DRV35_IFDET_BLUE_LED = DRV_IFDET_BLUE_LED_EN[35]? BLUE_DAT[35] : 1'bz;

endmodule